module half_adder(S,C,x,y);
    output S,C;
    input x,y;
    
    xor (S,x,y);
    and (C,x,y);
endmodule
